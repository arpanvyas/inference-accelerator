../../reg_intf/hdl/interface_regfile.sv