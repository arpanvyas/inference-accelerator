../../convolver/hdl/fifo_memory.sv