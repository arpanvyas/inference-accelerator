../../pool_nl/rtl/line_buffer_pool.sv