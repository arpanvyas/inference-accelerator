../../reg_intf/hdl/regfile_pool.sv