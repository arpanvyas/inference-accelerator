module register_top(

);
