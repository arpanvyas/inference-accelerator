../../top/rtl/controller.sv