../../reg_intf/hdl/regfile_nl.sv