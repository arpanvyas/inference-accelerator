../../pe_array/hdl/dense_latch.sv