../../convolver/hdl/shift_register9.sv