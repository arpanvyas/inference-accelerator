../../top/rtl/inference_accelerator.sv