`include "header.vh"
module host_system(
    input rst,
    input clk,
    input [1:0] input_bus1_PE,
    input [1:0] input_2_PE,
    output[1:0] output_1_PE
    );





endmodule
