../../top/header/header.vh