../../memory_bank/hdl/memory_buffer.sv