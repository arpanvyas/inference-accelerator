../../convolver/hdl/shift_register3.sv