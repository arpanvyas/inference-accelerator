../../reg_intf/hdl/regfile_fc.sv