../../reg_intf/hdl/reg_intf.sv