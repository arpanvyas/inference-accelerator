../../convolver/hdl/filter_buffer.sv