../../top/rtl/dense.sv