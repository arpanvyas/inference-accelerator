../../pool_nl/rtl/pooling.sv