../../convolver/hdl/line_fifo.sv