../../top/rtl/external_memory.sv