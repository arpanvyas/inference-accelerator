../../top/rtl/program_driver.sv