../../memory_bank/hdl/interface_buffer.sv