/home/vonfaust/data/accelerator/design/modules/top/rtl/buffer_pea_mux.sv