../../top/rtl/interface_extmem.sv