../../reg_intf/hdl/reg_intf_mux.sv