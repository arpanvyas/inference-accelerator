../../convolver/hdl/line_buffer.sv