../../reg_intf/hdl/spi_slave.sv