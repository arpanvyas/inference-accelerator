../../convolver/hdl/mac.sv