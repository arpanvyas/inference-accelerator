../../top/rtl/host.sv