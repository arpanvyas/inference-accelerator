../../pe_array/hdl/interface_pe_array.sv