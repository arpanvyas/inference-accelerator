../../top/header/user_tasks.vh