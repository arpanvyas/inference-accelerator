interface interface_extmem;

logic   we;
logic   re;
logic   [23:0]      rd_addr;
logic   [23:0]      wr_addr;
logic   [31:0]      rd_data;
logic   [31:0]      wr_data;

endinterface;
