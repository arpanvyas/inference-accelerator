../../pool_nl/rtl/adder_tree.sv