../../pe_array/hdl/PE_array.sv