../../pool_nl/rtl/densing.sv