../../reg_intf/hdl/regfile_general.sv