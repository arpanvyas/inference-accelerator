/home/vonfaust/data/accelerator/design/modules/top/rtl/computation_controller.sv