../../pool_nl/rtl/non_linearity.sv