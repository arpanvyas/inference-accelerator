interface intf();

logic   clk;
logic   rst;

logic   SCLK;
logic   SS;
logic   MOSI;
logic   MISO;

endinterface
