../../reg_intf/hdl/regfile_dense.sv