../../top/rtl/program_memory.sv