../../memory_bank/hdl/memory_bank.sv