../../reg_intf/hdl/register_top.sv