../../convolver/hdl/convolver.sv