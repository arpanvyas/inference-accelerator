../../convolver/hdl/shift_register2.sv