`ifndef SPI_HEADER
`define SPI_HEADER


`define NUM_SLAVES 1
`define PKT_SIZE  32



`endif
