../../top/rtl/pool.sv