task transaction;
    

endtask
