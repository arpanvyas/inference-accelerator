../../pe_array/hdl/PE.sv