../../convolver/hdl/multiplier.sv