../../top/rtl/conv.sv