../../reg_intf/hdl/sync_2s.sv