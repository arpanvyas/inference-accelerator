../../reg_intf/hdl/regfile_conv.sv